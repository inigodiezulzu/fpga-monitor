../../../../../../ip-core/monitor_1.0/hdl/monitor_control.vhd