../../../../../../ip-core/monitor_1.0/src/adc_manager.vhd