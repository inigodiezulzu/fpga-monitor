../../../../../../ip-core/monitor_1.0/src/spi_controller.vhd