../../../../../../ip-core/monitor_1.0/src/edge_detector.vhd