../../../../../../ip-core/monitor_1.0/src/counter.vhd