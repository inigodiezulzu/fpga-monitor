../../../../../../ip-core/monitor_1.0/src/bram_dualport.vhd