../../../../../../ip-core/monitor_1.0/src/fifo.vhd