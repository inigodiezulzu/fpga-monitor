../../../../../../ip-core/monitor_1.0/src/probes_trigger_module.vhd