../../../../../../ip-core/monitor_1.0/hdl/monitor_v1_0.vhd