../../../../../../ip-core/monitor_1.0/src/events_detector.vhd